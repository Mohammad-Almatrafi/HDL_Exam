// module multiplier (
//     input  [3:0] a,
//     input  [3:0] b,
//     output [7:0] y
// );


// nbitAdder #(.n(4))(.a(),.b(),.cin(),.y(),.cOut());




// endmodule
